// Timescale 
`timescale 1ns/1ps 
// Include source files 
`include "ips/pkgs/top_pkg.sv"
`include "ips/pkgs/prim_util_pkg.sv"
`include "ips/pkgs/prim_mubi_pkg.sv"
`include "ips/pkgs/prim_secded_pkg.sv"
`include "ips/pkgs/tlul_pkg.sv"
`include "tb/tlul_utils.sv"
`include "tb/tlul_if.sv"
`include "rtl/spi_host_reg_pkg.sv"
`ifndef SYN
  `include "rtl/spi_host.v"
`else
  `include "verilog/primitives.v"
  `include "verilog/sky130_fd_sc_hd.v"
  `include "syn/spi_host_synth.v"
`endif
