module twiddle_rom #(
  parameter int N = 1024,
  parameter int WIDTH = 16
)(
  input  logic [8:0] addr,
  output logic signed [WIDTH-1:0] re,
  output logic signed [WIDTH-1:0] im
);

  // ROM arrays to hold precomputed twiddle factors
  logic signed [WIDTH-1:0] rom_re [0:N/2-1];
  logic signed [WIDTH-1:0] rom_im [0:N/2-1];

  initial begin
    rom_re[0] = 32768;
    rom_re[1] = 32767;
    rom_re[2] = 32766;
    rom_re[3] = 32762;
    rom_re[4] = 32758;
    rom_re[5] = 32753;
    rom_re[6] = 32746;
    rom_re[7] = 32738;
    rom_re[8] = 32729;
    rom_re[9] = 32718;
    rom_re[10] = 32706;
    rom_re[11] = 32693;
    rom_re[12] = 32679;
    rom_re[13] = 32664;
    rom_re[14] = 32647;
    rom_re[15] = 32629;
    rom_re[16] = 32610;
    rom_re[17] = 32590;
    rom_re[18] = 32568;
    rom_re[19] = 32546;
    rom_re[20] = 32522;
    rom_re[21] = 32496;
    rom_re[22] = 32470;
    rom_re[23] = 32442;
    rom_re[24] = 32413;
    rom_re[25] = 32383;
    rom_re[26] = 32352;
    rom_re[27] = 32319;
    rom_re[28] = 32286;
    rom_re[29] = 32251;
    rom_re[30] = 32214;
    rom_re[31] = 32177;
    rom_re[32] = 32138;
    rom_re[33] = 32099;
    rom_re[34] = 32058;
    rom_re[35] = 32015;
    rom_re[36] = 31972;
    rom_re[37] = 31927;
    rom_re[38] = 31881;
    rom_re[39] = 31834;
    rom_re[40] = 31786;
    rom_re[41] = 31737;
    rom_re[42] = 31686;
    rom_re[43] = 31634;
    rom_re[44] = 31581;
    rom_re[45] = 31527;
    rom_re[46] = 31471;
    rom_re[47] = 31415;
    rom_re[48] = 31357;
    rom_re[49] = 31298;
    rom_re[50] = 31238;
    rom_re[51] = 31177;
    rom_re[52] = 31114;
    rom_re[53] = 31050;
    rom_re[54] = 30986;
    rom_re[55] = 30920;
    rom_re[56] = 30853;
    rom_re[57] = 30784;
    rom_re[58] = 30715;
    rom_re[59] = 30644;
    rom_re[60] = 30572;
    rom_re[61] = 30499;
    rom_re[62] = 30425;
    rom_re[63] = 30350;
    rom_re[64] = 30274;
    rom_re[65] = 30196;
    rom_re[66] = 30118;
    rom_re[67] = 30038;
    rom_re[68] = 29957;
    rom_re[69] = 29875;
    rom_re[70] = 29792;
    rom_re[71] = 29707;
    rom_re[72] = 29622;
    rom_re[73] = 29535;
    rom_re[74] = 29448;
    rom_re[75] = 29359;
    rom_re[76] = 29269;
    rom_re[77] = 29178;
    rom_re[78] = 29086;
    rom_re[79] = 28993;
    rom_re[80] = 28899;
    rom_re[81] = 28803;
    rom_re[82] = 28707;
    rom_re[83] = 28610;
    rom_re[84] = 28511;
    rom_re[85] = 28411;
    rom_re[86] = 28311;
    rom_re[87] = 28209;
    rom_re[88] = 28106;
    rom_re[89] = 28002;
    rom_re[90] = 27897;
    rom_re[91] = 27791;
    rom_re[92] = 27684;
    rom_re[93] = 27576;
    rom_re[94] = 27467;
    rom_re[95] = 27357;
    rom_re[96] = 27246;
    rom_re[97] = 27133;
    rom_re[98] = 27020;
    rom_re[99] = 26906;
    rom_re[100] = 26791;
    rom_re[101] = 26674;
    rom_re[102] = 26557;
    rom_re[103] = 26439;
    rom_re[104] = 26320;
    rom_re[105] = 26199;
    rom_re[106] = 26078;
    rom_re[107] = 25956;
    rom_re[108] = 25833;
    rom_re[109] = 25708;
    rom_re[110] = 25583;
    rom_re[111] = 25457;
    rom_re[112] = 25330;
    rom_re[113] = 25202;
    rom_re[114] = 25073;
    rom_re[115] = 24943;
    rom_re[116] = 24812;
    rom_re[117] = 24680;
    rom_re[118] = 24548;
    rom_re[119] = 24414;
    rom_re[120] = 24279;
    rom_re[121] = 24144;
    rom_re[122] = 24008;
    rom_re[123] = 23870;
    rom_re[124] = 23732;
    rom_re[125] = 23593;
    rom_re[126] = 23453;
    rom_re[127] = 23312;
    rom_re[128] = 23170;
    rom_re[129] = 23028;
    rom_re[130] = 22884;
    rom_re[131] = 22740;
    rom_re[132] = 22595;
    rom_re[133] = 22449;
    rom_re[134] = 22302;
    rom_re[135] = 22154;
    rom_re[136] = 22006;
    rom_re[137] = 21856;
    rom_re[138] = 21706;
    rom_re[139] = 21555;
    rom_re[140] = 21403;
    rom_re[141] = 21251;
    rom_re[142] = 21097;
    rom_re[143] = 20943;
    rom_re[144] = 20788;
    rom_re[145] = 20632;
    rom_re[146] = 20475;
    rom_re[147] = 20318;
    rom_re[148] = 20160;
    rom_re[149] = 20001;
    rom_re[150] = 19841;
    rom_re[151] = 19681;
    rom_re[152] = 19520;
    rom_re[153] = 19358;
    rom_re[154] = 19195;
    rom_re[155] = 19032;
    rom_re[156] = 18868;
    rom_re[157] = 18703;
    rom_re[158] = 18538;
    rom_re[159] = 18372;
    rom_re[160] = 18205;
    rom_re[161] = 18037;
    rom_re[162] = 17869;
    rom_re[163] = 17700;
    rom_re[164] = 17531;
    rom_re[165] = 17361;
    rom_re[166] = 17190;
    rom_re[167] = 17018;
    rom_re[168] = 16846;
    rom_re[169] = 16673;
    rom_re[170] = 16500;
    rom_re[171] = 16326;
    rom_re[172] = 16151;
    rom_re[173] = 15976;
    rom_re[174] = 15800;
    rom_re[175] = 15624;
    rom_re[176] = 15447;
    rom_re[177] = 15269;
    rom_re[178] = 15091;
    rom_re[179] = 14912;
    rom_re[180] = 14733;
    rom_re[181] = 14553;
    rom_re[182] = 14373;
    rom_re[183] = 14192;
    rom_re[184] = 14010;
    rom_re[185] = 13828;
    rom_re[186] = 13646;
    rom_re[187] = 13463;
    rom_re[188] = 13279;
    rom_re[189] = 13095;
    rom_re[190] = 12910;
    rom_re[191] = 12725;
    rom_re[192] = 12540;
    rom_re[193] = 12354;
    rom_re[194] = 12167;
    rom_re[195] = 11980;
    rom_re[196] = 11793;
    rom_re[197] = 11605;
    rom_re[198] = 11417;
    rom_re[199] = 11228;
    rom_re[200] = 11039;
    rom_re[201] = 10850;
    rom_re[202] = 10660;
    rom_re[203] = 10469;
    rom_re[204] = 10279;
    rom_re[205] = 10088;
    rom_re[206] = 9896;
    rom_re[207] = 9704;
    rom_re[208] = 9512;
    rom_re[209] = 9319;
    rom_re[210] = 9127;
    rom_re[211] = 8933;
    rom_re[212] = 8740;
    rom_re[213] = 8546;
    rom_re[214] = 8351;
    rom_re[215] = 8157;
    rom_re[216] = 7962;
    rom_re[217] = 7767;
    rom_re[218] = 7571;
    rom_re[219] = 7376;
    rom_re[220] = 7180;
    rom_re[221] = 6983;
    rom_re[222] = 6787;
    rom_re[223] = 6590;
    rom_re[224] = 6393;
    rom_re[225] = 6195;
    rom_re[226] = 5998;
    rom_re[227] = 5800;
    rom_re[228] = 5602;
    rom_re[229] = 5404;
    rom_re[230] = 5205;
    rom_re[231] = 5007;
    rom_re[232] = 4808;
    rom_re[233] = 4609;
    rom_re[234] = 4410;
    rom_re[235] = 4211;
    rom_re[236] = 4011;
    rom_re[237] = 3812;
    rom_re[238] = 3612;
    rom_re[239] = 3412;
    rom_re[240] = 3212;
    rom_re[241] = 3012;
    rom_re[242] = 2811;
    rom_re[243] = 2611;
    rom_re[244] = 2411;
    rom_re[245] = 2210;
    rom_re[246] = 2009;
    rom_re[247] = 1809;
    rom_re[248] = 1608;
    rom_re[249] = 1407;
    rom_re[250] = 1206;
    rom_re[251] = 1005;
    rom_re[252] = 804;
    rom_re[253] = 603;
    rom_re[254] = 402;
    rom_re[255] = 201;
    rom_re[256] = 0;
    rom_re[257] = -201;
    rom_re[258] = -402;
    rom_re[259] = -603;
    rom_re[260] = -804;
    rom_re[261] = -1005;
    rom_re[262] = -1206;
    rom_re[263] = -1407;
    rom_re[264] = -1608;
    rom_re[265] = -1809;
    rom_re[266] = -2009;
    rom_re[267] = -2210;
    rom_re[268] = -2411;
    rom_re[269] = -2611;
    rom_re[270] = -2811;
    rom_re[271] = -3012;
    rom_re[272] = -3212;
    rom_re[273] = -3412;
    rom_re[274] = -3612;
    rom_re[275] = -3812;
    rom_re[276] = -4011;
    rom_re[277] = -4211;
    rom_re[278] = -4410;
    rom_re[279] = -4609;
    rom_re[280] = -4808;
    rom_re[281] = -5007;
    rom_re[282] = -5205;
    rom_re[283] = -5404;
    rom_re[284] = -5602;
    rom_re[285] = -5800;
    rom_re[286] = -5998;
    rom_re[287] = -6195;
    rom_re[288] = -6393;
    rom_re[289] = -6590;
    rom_re[290] = -6787;
    rom_re[291] = -6983;
    rom_re[292] = -7180;
    rom_re[293] = -7376;
    rom_re[294] = -7571;
    rom_re[295] = -7767;
    rom_re[296] = -7962;
    rom_re[297] = -8157;
    rom_re[298] = -8351;
    rom_re[299] = -8546;
    rom_re[300] = -8740;
    rom_re[301] = -8933;
    rom_re[302] = -9127;
    rom_re[303] = -9319;
    rom_re[304] = -9512;
    rom_re[305] = -9704;
    rom_re[306] = -9896;
    rom_re[307] = -10088;
    rom_re[308] = -10279;
    rom_re[309] = -10469;
    rom_re[310] = -10660;
    rom_re[311] = -10850;
    rom_re[312] = -11039;
    rom_re[313] = -11228;
    rom_re[314] = -11417;
    rom_re[315] = -11605;
    rom_re[316] = -11793;
    rom_re[317] = -11980;
    rom_re[318] = -12167;
    rom_re[319] = -12354;
    rom_re[320] = -12540;
    rom_re[321] = -12725;
    rom_re[322] = -12910;
    rom_re[323] = -13095;
    rom_re[324] = -13279;
    rom_re[325] = -13463;
    rom_re[326] = -13646;
    rom_re[327] = -13828;
    rom_re[328] = -14010;
    rom_re[329] = -14192;
    rom_re[330] = -14373;
    rom_re[331] = -14553;
    rom_re[332] = -14733;
    rom_re[333] = -14912;
    rom_re[334] = -15091;
    rom_re[335] = -15269;
    rom_re[336] = -15447;
    rom_re[337] = -15624;
    rom_re[338] = -15800;
    rom_re[339] = -15976;
    rom_re[340] = -16151;
    rom_re[341] = -16326;
    rom_re[342] = -16500;
    rom_re[343] = -16673;
    rom_re[344] = -16846;
    rom_re[345] = -17018;
    rom_re[346] = -17190;
    rom_re[347] = -17361;
    rom_re[348] = -17531;
    rom_re[349] = -17700;
    rom_re[350] = -17869;
    rom_re[351] = -18037;
    rom_re[352] = -18205;
    rom_re[353] = -18372;
    rom_re[354] = -18538;
    rom_re[355] = -18703;
    rom_re[356] = -18868;
    rom_re[357] = -19032;
    rom_re[358] = -19195;
    rom_re[359] = -19358;
    rom_re[360] = -19520;
    rom_re[361] = -19681;
    rom_re[362] = -19841;
    rom_re[363] = -20001;
    rom_re[364] = -20160;
    rom_re[365] = -20318;
    rom_re[366] = -20475;
    rom_re[367] = -20632;
    rom_re[368] = -20788;
    rom_re[369] = -20943;
    rom_re[370] = -21097;
    rom_re[371] = -21251;
    rom_re[372] = -21403;
    rom_re[373] = -21555;
    rom_re[374] = -21706;
    rom_re[375] = -21856;
    rom_re[376] = -22006;
    rom_re[377] = -22154;
    rom_re[378] = -22302;
    rom_re[379] = -22449;
    rom_re[380] = -22595;
    rom_re[381] = -22740;
    rom_re[382] = -22884;
    rom_re[383] = -23028;
    rom_re[384] = -23170;
    rom_re[385] = -23312;
    rom_re[386] = -23453;
    rom_re[387] = -23593;
    rom_re[388] = -23732;
    rom_re[389] = -23870;
    rom_re[390] = -24008;
    rom_re[391] = -24144;
    rom_re[392] = -24279;
    rom_re[393] = -24414;
    rom_re[394] = -24548;
    rom_re[395] = -24680;
    rom_re[396] = -24812;
    rom_re[397] = -24943;
    rom_re[398] = -25073;
    rom_re[399] = -25202;
    rom_re[400] = -25330;
    rom_re[401] = -25457;
    rom_re[402] = -25583;
    rom_re[403] = -25708;
    rom_re[404] = -25833;
    rom_re[405] = -25956;
    rom_re[406] = -26078;
    rom_re[407] = -26199;
    rom_re[408] = -26320;
    rom_re[409] = -26439;
    rom_re[410] = -26557;
    rom_re[411] = -26674;
    rom_re[412] = -26791;
    rom_re[413] = -26906;
    rom_re[414] = -27020;
    rom_re[415] = -27133;
    rom_re[416] = -27246;
    rom_re[417] = -27357;
    rom_re[418] = -27467;
    rom_re[419] = -27576;
    rom_re[420] = -27684;
    rom_re[421] = -27791;
    rom_re[422] = -27897;
    rom_re[423] = -28002;
    rom_re[424] = -28106;
    rom_re[425] = -28209;
    rom_re[426] = -28311;
    rom_re[427] = -28411;
    rom_re[428] = -28511;
    rom_re[429] = -28610;
    rom_re[430] = -28707;
    rom_re[431] = -28803;
    rom_re[432] = -28899;
    rom_re[433] = -28993;
    rom_re[434] = -29086;
    rom_re[435] = -29178;
    rom_re[436] = -29269;
    rom_re[437] = -29359;
    rom_re[438] = -29448;
    rom_re[439] = -29535;
    rom_re[440] = -29622;
    rom_re[441] = -29707;
    rom_re[442] = -29792;
    rom_re[443] = -29875;
    rom_re[444] = -29957;
    rom_re[445] = -30038;
    rom_re[446] = -30118;
    rom_re[447] = -30196;
    rom_re[448] = -30274;
    rom_re[449] = -30350;
    rom_re[450] = -30425;
    rom_re[451] = -30499;
    rom_re[452] = -30572;
    rom_re[453] = -30644;
    rom_re[454] = -30715;
    rom_re[455] = -30784;
    rom_re[456] = -30853;
    rom_re[457] = -30920;
    rom_re[458] = -30986;
    rom_re[459] = -31050;
    rom_re[460] = -31114;
    rom_re[461] = -31177;
    rom_re[462] = -31238;
    rom_re[463] = -31298;
    rom_re[464] = -31357;
    rom_re[465] = -31415;
    rom_re[466] = -31471;
    rom_re[467] = -31527;
    rom_re[468] = -31581;
    rom_re[469] = -31634;
    rom_re[470] = -31686;
    rom_re[471] = -31737;
    rom_re[472] = -31786;
    rom_re[473] = -31834;
    rom_re[474] = -31881;
    rom_re[475] = -31927;
    rom_re[476] = -31972;
    rom_re[477] = -32015;
    rom_re[478] = -32058;
    rom_re[479] = -32099;
    rom_re[480] = -32138;
    rom_re[481] = -32177;
    rom_re[482] = -32214;
    rom_re[483] = -32251;
    rom_re[484] = -32286;
    rom_re[485] = -32319;
    rom_re[486] = -32352;
    rom_re[487] = -32383;
    rom_re[488] = -32413;
    rom_re[489] = -32442;
    rom_re[490] = -32470;
    rom_re[491] = -32496;
    rom_re[492] = -32522;
    rom_re[493] = -32546;
    rom_re[494] = -32568;
    rom_re[495] = -32590;
    rom_re[496] = -32610;
    rom_re[497] = -32629;
    rom_re[498] = -32647;
    rom_re[499] = -32664;
    rom_re[500] = -32679;
    rom_re[501] = -32693;
    rom_re[502] = -32706;
    rom_re[503] = -32718;
    rom_re[504] = -32729;
    rom_re[505] = -32738;
    rom_re[506] = -32746;
    rom_re[507] = -32753;
    rom_re[508] = -32758;
    rom_re[509] = -32762;
    rom_re[510] = -32766;
    rom_re[511] = -32767;
    rom_im[0] = 0;
    rom_im[1] = -201;
    rom_im[2] = -402;
    rom_im[3] = -603;
    rom_im[4] = -804;
    rom_im[5] = -1005;
    rom_im[6] = -1206;
    rom_im[7] = -1407;
    rom_im[8] = -1608;
    rom_im[9] = -1809;
    rom_im[10] = -2009;
    rom_im[11] = -2210;
    rom_im[12] = -2411;
    rom_im[13] = -2611;
    rom_im[14] = -2811;
    rom_im[15] = -3012;
    rom_im[16] = -3212;
    rom_im[17] = -3412;
    rom_im[18] = -3612;
    rom_im[19] = -3812;
    rom_im[20] = -4011;
    rom_im[21] = -4211;
    rom_im[22] = -4410;
    rom_im[23] = -4609;
    rom_im[24] = -4808;
    rom_im[25] = -5007;
    rom_im[26] = -5205;
    rom_im[27] = -5404;
    rom_im[28] = -5602;
    rom_im[29] = -5800;
    rom_im[30] = -5998;
    rom_im[31] = -6195;
    rom_im[32] = -6393;
    rom_im[33] = -6590;
    rom_im[34] = -6787;
    rom_im[35] = -6983;
    rom_im[36] = -7180;
    rom_im[37] = -7376;
    rom_im[38] = -7571;
    rom_im[39] = -7767;
    rom_im[40] = -7962;
    rom_im[41] = -8157;
    rom_im[42] = -8351;
    rom_im[43] = -8546;
    rom_im[44] = -8740;
    rom_im[45] = -8933;
    rom_im[46] = -9127;
    rom_im[47] = -9319;
    rom_im[48] = -9512;
    rom_im[49] = -9704;
    rom_im[50] = -9896;
    rom_im[51] = -10088;
    rom_im[52] = -10279;
    rom_im[53] = -10469;
    rom_im[54] = -10660;
    rom_im[55] = -10850;
    rom_im[56] = -11039;
    rom_im[57] = -11228;
    rom_im[58] = -11417;
    rom_im[59] = -11605;
    rom_im[60] = -11793;
    rom_im[61] = -11980;
    rom_im[62] = -12167;
    rom_im[63] = -12354;
    rom_im[64] = -12540;
    rom_im[65] = -12725;
    rom_im[66] = -12910;
    rom_im[67] = -13095;
    rom_im[68] = -13279;
    rom_im[69] = -13463;
    rom_im[70] = -13646;
    rom_im[71] = -13828;
    rom_im[72] = -14010;
    rom_im[73] = -14192;
    rom_im[74] = -14373;
    rom_im[75] = -14553;
    rom_im[76] = -14733;
    rom_im[77] = -14912;
    rom_im[78] = -15091;
    rom_im[79] = -15269;
    rom_im[80] = -15447;
    rom_im[81] = -15624;
    rom_im[82] = -15800;
    rom_im[83] = -15976;
    rom_im[84] = -16151;
    rom_im[85] = -16326;
    rom_im[86] = -16500;
    rom_im[87] = -16673;
    rom_im[88] = -16846;
    rom_im[89] = -17018;
    rom_im[90] = -17190;
    rom_im[91] = -17361;
    rom_im[92] = -17531;
    rom_im[93] = -17700;
    rom_im[94] = -17869;
    rom_im[95] = -18037;
    rom_im[96] = -18205;
    rom_im[97] = -18372;
    rom_im[98] = -18538;
    rom_im[99] = -18703;
    rom_im[100] = -18868;
    rom_im[101] = -19032;
    rom_im[102] = -19195;
    rom_im[103] = -19358;
    rom_im[104] = -19520;
    rom_im[105] = -19681;
    rom_im[106] = -19841;
    rom_im[107] = -20001;
    rom_im[108] = -20160;
    rom_im[109] = -20318;
    rom_im[110] = -20475;
    rom_im[111] = -20632;
    rom_im[112] = -20788;
    rom_im[113] = -20943;
    rom_im[114] = -21097;
    rom_im[115] = -21251;
    rom_im[116] = -21403;
    rom_im[117] = -21555;
    rom_im[118] = -21706;
    rom_im[119] = -21856;
    rom_im[120] = -22006;
    rom_im[121] = -22154;
    rom_im[122] = -22302;
    rom_im[123] = -22449;
    rom_im[124] = -22595;
    rom_im[125] = -22740;
    rom_im[126] = -22884;
    rom_im[127] = -23028;
    rom_im[128] = -23170;
    rom_im[129] = -23312;
    rom_im[130] = -23453;
    rom_im[131] = -23593;
    rom_im[132] = -23732;
    rom_im[133] = -23870;
    rom_im[134] = -24008;
    rom_im[135] = -24144;
    rom_im[136] = -24279;
    rom_im[137] = -24414;
    rom_im[138] = -24548;
    rom_im[139] = -24680;
    rom_im[140] = -24812;
    rom_im[141] = -24943;
    rom_im[142] = -25073;
    rom_im[143] = -25202;
    rom_im[144] = -25330;
    rom_im[145] = -25457;
    rom_im[146] = -25583;
    rom_im[147] = -25708;
    rom_im[148] = -25833;
    rom_im[149] = -25956;
    rom_im[150] = -26078;
    rom_im[151] = -26199;
    rom_im[152] = -26320;
    rom_im[153] = -26439;
    rom_im[154] = -26557;
    rom_im[155] = -26674;
    rom_im[156] = -26791;
    rom_im[157] = -26906;
    rom_im[158] = -27020;
    rom_im[159] = -27133;
    rom_im[160] = -27246;
    rom_im[161] = -27357;
    rom_im[162] = -27467;
    rom_im[163] = -27576;
    rom_im[164] = -27684;
    rom_im[165] = -27791;
    rom_im[166] = -27897;
    rom_im[167] = -28002;
    rom_im[168] = -28106;
    rom_im[169] = -28209;
    rom_im[170] = -28311;
    rom_im[171] = -28411;
    rom_im[172] = -28511;
    rom_im[173] = -28610;
    rom_im[174] = -28707;
    rom_im[175] = -28803;
    rom_im[176] = -28899;
    rom_im[177] = -28993;
    rom_im[178] = -29086;
    rom_im[179] = -29178;
    rom_im[180] = -29269;
    rom_im[181] = -29359;
    rom_im[182] = -29448;
    rom_im[183] = -29535;
    rom_im[184] = -29622;
    rom_im[185] = -29707;
    rom_im[186] = -29792;
    rom_im[187] = -29875;
    rom_im[188] = -29957;
    rom_im[189] = -30038;
    rom_im[190] = -30118;
    rom_im[191] = -30196;
    rom_im[192] = -30274;
    rom_im[193] = -30350;
    rom_im[194] = -30425;
    rom_im[195] = -30499;
    rom_im[196] = -30572;
    rom_im[197] = -30644;
    rom_im[198] = -30715;
    rom_im[199] = -30784;
    rom_im[200] = -30853;
    rom_im[201] = -30920;
    rom_im[202] = -30986;
    rom_im[203] = -31050;
    rom_im[204] = -31114;
    rom_im[205] = -31177;
    rom_im[206] = -31238;
    rom_im[207] = -31298;
    rom_im[208] = -31357;
    rom_im[209] = -31415;
    rom_im[210] = -31471;
    rom_im[211] = -31527;
    rom_im[212] = -31581;
    rom_im[213] = -31634;
    rom_im[214] = -31686;
    rom_im[215] = -31737;
    rom_im[216] = -31786;
    rom_im[217] = -31834;
    rom_im[218] = -31881;
    rom_im[219] = -31927;
    rom_im[220] = -31972;
    rom_im[221] = -32015;
    rom_im[222] = -32058;
    rom_im[223] = -32099;
    rom_im[224] = -32138;
    rom_im[225] = -32177;
    rom_im[226] = -32214;
    rom_im[227] = -32251;
    rom_im[228] = -32286;
    rom_im[229] = -32319;
    rom_im[230] = -32352;
    rom_im[231] = -32383;
    rom_im[232] = -32413;
    rom_im[233] = -32442;
    rom_im[234] = -32470;
    rom_im[235] = -32496;
    rom_im[236] = -32522;
    rom_im[237] = -32546;
    rom_im[238] = -32568;
    rom_im[239] = -32590;
    rom_im[240] = -32610;
    rom_im[241] = -32629;
    rom_im[242] = -32647;
    rom_im[243] = -32664;
    rom_im[244] = -32679;
    rom_im[245] = -32693;
    rom_im[246] = -32706;
    rom_im[247] = -32718;
    rom_im[248] = -32729;
    rom_im[249] = -32738;
    rom_im[250] = -32746;
    rom_im[251] = -32753;
    rom_im[252] = -32758;
    rom_im[253] = -32762;
    rom_im[254] = -32766;
    rom_im[255] = -32767;
    rom_im[256] = -32768;
    rom_im[257] = -32767;
    rom_im[258] = -32766;
    rom_im[259] = -32762;
    rom_im[260] = -32758;
    rom_im[261] = -32753;
    rom_im[262] = -32746;
    rom_im[263] = -32738;
    rom_im[264] = -32729;
    rom_im[265] = -32718;
    rom_im[266] = -32706;
    rom_im[267] = -32693;
    rom_im[268] = -32679;
    rom_im[269] = -32664;
    rom_im[270] = -32647;
    rom_im[271] = -32629;
    rom_im[272] = -32610;
    rom_im[273] = -32590;
    rom_im[274] = -32568;
    rom_im[275] = -32546;
    rom_im[276] = -32522;
    rom_im[277] = -32496;
    rom_im[278] = -32470;
    rom_im[279] = -32442;
    rom_im[280] = -32413;
    rom_im[281] = -32383;
    rom_im[282] = -32352;
    rom_im[283] = -32319;
    rom_im[284] = -32286;
    rom_im[285] = -32251;
    rom_im[286] = -32214;
    rom_im[287] = -32177;
    rom_im[288] = -32138;
    rom_im[289] = -32099;
    rom_im[290] = -32058;
    rom_im[291] = -32015;
    rom_im[292] = -31972;
    rom_im[293] = -31927;
    rom_im[294] = -31881;
    rom_im[295] = -31834;
    rom_im[296] = -31786;
    rom_im[297] = -31737;
    rom_im[298] = -31686;
    rom_im[299] = -31634;
    rom_im[300] = -31581;
    rom_im[301] = -31527;
    rom_im[302] = -31471;
    rom_im[303] = -31415;
    rom_im[304] = -31357;
    rom_im[305] = -31298;
    rom_im[306] = -31238;
    rom_im[307] = -31177;
    rom_im[308] = -31114;
    rom_im[309] = -31050;
    rom_im[310] = -30986;
    rom_im[311] = -30920;
    rom_im[312] = -30853;
    rom_im[313] = -30784;
    rom_im[314] = -30715;
    rom_im[315] = -30644;
    rom_im[316] = -30572;
    rom_im[317] = -30499;
    rom_im[318] = -30425;
    rom_im[319] = -30350;
    rom_im[320] = -30274;
    rom_im[321] = -30196;
    rom_im[322] = -30118;
    rom_im[323] = -30038;
    rom_im[324] = -29957;
    rom_im[325] = -29875;
    rom_im[326] = -29792;
    rom_im[327] = -29707;
    rom_im[328] = -29622;
    rom_im[329] = -29535;
    rom_im[330] = -29448;
    rom_im[331] = -29359;
    rom_im[332] = -29269;
    rom_im[333] = -29178;
    rom_im[334] = -29086;
    rom_im[335] = -28993;
    rom_im[336] = -28899;
    rom_im[337] = -28803;
    rom_im[338] = -28707;
    rom_im[339] = -28610;
    rom_im[340] = -28511;
    rom_im[341] = -28411;
    rom_im[342] = -28311;
    rom_im[343] = -28209;
    rom_im[344] = -28106;
    rom_im[345] = -28002;
    rom_im[346] = -27897;
    rom_im[347] = -27791;
    rom_im[348] = -27684;
    rom_im[349] = -27576;
    rom_im[350] = -27467;
    rom_im[351] = -27357;
    rom_im[352] = -27246;
    rom_im[353] = -27133;
    rom_im[354] = -27020;
    rom_im[355] = -26906;
    rom_im[356] = -26791;
    rom_im[357] = -26674;
    rom_im[358] = -26557;
    rom_im[359] = -26439;
    rom_im[360] = -26320;
    rom_im[361] = -26199;
    rom_im[362] = -26078;
    rom_im[363] = -25956;
    rom_im[364] = -25833;
    rom_im[365] = -25708;
    rom_im[366] = -25583;
    rom_im[367] = -25457;
    rom_im[368] = -25330;
    rom_im[369] = -25202;
    rom_im[370] = -25073;
    rom_im[371] = -24943;
    rom_im[372] = -24812;
    rom_im[373] = -24680;
    rom_im[374] = -24548;
    rom_im[375] = -24414;
    rom_im[376] = -24279;
    rom_im[377] = -24144;
    rom_im[378] = -24008;
    rom_im[379] = -23870;
    rom_im[380] = -23732;
    rom_im[381] = -23593;
    rom_im[382] = -23453;
    rom_im[383] = -23312;
    rom_im[384] = -23170;
    rom_im[385] = -23028;
    rom_im[386] = -22884;
    rom_im[387] = -22740;
    rom_im[388] = -22595;
    rom_im[389] = -22449;
    rom_im[390] = -22302;
    rom_im[391] = -22154;
    rom_im[392] = -22006;
    rom_im[393] = -21856;
    rom_im[394] = -21706;
    rom_im[395] = -21555;
    rom_im[396] = -21403;
    rom_im[397] = -21251;
    rom_im[398] = -21097;
    rom_im[399] = -20943;
    rom_im[400] = -20788;
    rom_im[401] = -20632;
    rom_im[402] = -20475;
    rom_im[403] = -20318;
    rom_im[404] = -20160;
    rom_im[405] = -20001;
    rom_im[406] = -19841;
    rom_im[407] = -19681;
    rom_im[408] = -19520;
    rom_im[409] = -19358;
    rom_im[410] = -19195;
    rom_im[411] = -19032;
    rom_im[412] = -18868;
    rom_im[413] = -18703;
    rom_im[414] = -18538;
    rom_im[415] = -18372;
    rom_im[416] = -18205;
    rom_im[417] = -18037;
    rom_im[418] = -17869;
    rom_im[419] = -17700;
    rom_im[420] = -17531;
    rom_im[421] = -17361;
    rom_im[422] = -17190;
    rom_im[423] = -17018;
    rom_im[424] = -16846;
    rom_im[425] = -16673;
    rom_im[426] = -16500;
    rom_im[427] = -16326;
    rom_im[428] = -16151;
    rom_im[429] = -15976;
    rom_im[430] = -15800;
    rom_im[431] = -15624;
    rom_im[432] = -15447;
    rom_im[433] = -15269;
    rom_im[434] = -15091;
    rom_im[435] = -14912;
    rom_im[436] = -14733;
    rom_im[437] = -14553;
    rom_im[438] = -14373;
    rom_im[439] = -14192;
    rom_im[440] = -14010;
    rom_im[441] = -13828;
    rom_im[442] = -13646;
    rom_im[443] = -13463;
    rom_im[444] = -13279;
    rom_im[445] = -13095;
    rom_im[446] = -12910;
    rom_im[447] = -12725;
    rom_im[448] = -12540;
    rom_im[449] = -12354;
    rom_im[450] = -12167;
    rom_im[451] = -11980;
    rom_im[452] = -11793;
    rom_im[453] = -11605;
    rom_im[454] = -11417;
    rom_im[455] = -11228;
    rom_im[456] = -11039;
    rom_im[457] = -10850;
    rom_im[458] = -10660;
    rom_im[459] = -10469;
    rom_im[460] = -10279;
    rom_im[461] = -10088;
    rom_im[462] = -9896;
    rom_im[463] = -9704;
    rom_im[464] = -9512;
    rom_im[465] = -9319;
    rom_im[466] = -9127;
    rom_im[467] = -8933;
    rom_im[468] = -8740;
    rom_im[469] = -8546;
    rom_im[470] = -8351;
    rom_im[471] = -8157;
    rom_im[472] = -7962;
    rom_im[473] = -7767;
    rom_im[474] = -7571;
    rom_im[475] = -7376;
    rom_im[476] = -7180;
    rom_im[477] = -6983;
    rom_im[478] = -6787;
    rom_im[479] = -6590;
    rom_im[480] = -6393;
    rom_im[481] = -6195;
    rom_im[482] = -5998;
    rom_im[483] = -5800;
    rom_im[484] = -5602;
    rom_im[485] = -5404;
    rom_im[486] = -5205;
    rom_im[487] = -5007;
    rom_im[488] = -4808;
    rom_im[489] = -4609;
    rom_im[490] = -4410;
    rom_im[491] = -4211;
    rom_im[492] = -4011;
    rom_im[493] = -3812;
    rom_im[494] = -3612;
    rom_im[495] = -3412;
    rom_im[496] = -3212;
    rom_im[497] = -3012;
    rom_im[498] = -2811;
    rom_im[499] = -2611;
    rom_im[500] = -2411;
    rom_im[501] = -2210;
    rom_im[502] = -2009;
    rom_im[503] = -1809;
    rom_im[504] = -1608;
    rom_im[505] = -1407;
    rom_im[506] = -1206;
    rom_im[507] = -1005;
    rom_im[508] = -804;
    rom_im[509] = -603;
    rom_im[510] = -402;
    rom_im[511] = -201;
  end

  always_comb begin
    re = rom_re[addr];
    im = rom_im[addr];
  end

endmodule
