module twiddle_rom_256 #(
  parameter int N = 256,
  parameter int WIDTH = 16
)(
  input  logic [6:0] addr,
  output logic signed [WIDTH-1:0] re,
  output logic signed [WIDTH-1:0] im
);

  // ROM arrays to hold precomputed twiddle factors
  logic signed [WIDTH-1:0] rom_re [0:N/2-1];
  logic signed [WIDTH-1:0] rom_im [0:N/2-1];

  initial begin
    rom_re[0] = 32768;
    rom_re[1] = 32758;
    rom_re[2] = 32729;
    rom_re[3] = 32679;
    rom_re[4] = 32610;
    rom_re[5] = 32522;
    rom_re[6] = 32413;
    rom_re[7] = 32286;
    rom_re[8] = 32138;
    rom_re[9] = 31972;
    rom_re[10] = 31786;
    rom_re[11] = 31581;
    rom_re[12] = 31357;
    rom_re[13] = 31114;
    rom_re[14] = 30853;
    rom_re[15] = 30572;
    rom_re[16] = 30274;
    rom_re[17] = 29957;
    rom_re[18] = 29622;
    rom_re[19] = 29269;
    rom_re[20] = 28899;
    rom_re[21] = 28511;
    rom_re[22] = 28106;
    rom_re[23] = 27684;
    rom_re[24] = 27246;
    rom_re[25] = 26791;
    rom_re[26] = 26320;
    rom_re[27] = 25833;
    rom_re[28] = 25330;
    rom_re[29] = 24812;
    rom_re[30] = 24279;
    rom_re[31] = 23732;
    rom_re[32] = 23170;
    rom_re[33] = 22595;
    rom_re[34] = 22006;
    rom_re[35] = 21403;
    rom_re[36] = 20788;
    rom_re[37] = 20160;
    rom_re[38] = 19520;
    rom_re[39] = 18868;
    rom_re[40] = 18205;
    rom_re[41] = 17531;
    rom_re[42] = 16846;
    rom_re[43] = 16151;
    rom_re[44] = 15447;
    rom_re[45] = 14733;
    rom_re[46] = 14010;
    rom_re[47] = 13279;
    rom_re[48] = 12540;
    rom_re[49] = 11793;
    rom_re[50] = 11039;
    rom_re[51] = 10279;
    rom_re[52] = 9512;
    rom_re[53] = 8740;
    rom_re[54] = 7962;
    rom_re[55] = 7180;
    rom_re[56] = 6393;
    rom_re[57] = 5602;
    rom_re[58] = 4808;
    rom_re[59] = 4011;
    rom_re[60] = 3212;
    rom_re[61] = 2411;
    rom_re[62] = 1608;
    rom_re[63] = 804;
    rom_re[64] = 0;
    rom_re[65] = -804;
    rom_re[66] = -1608;
    rom_re[67] = -2411;
    rom_re[68] = -3212;
    rom_re[69] = -4011;
    rom_re[70] = -4808;
    rom_re[71] = -5602;
    rom_re[72] = -6393;
    rom_re[73] = -7180;
    rom_re[74] = -7962;
    rom_re[75] = -8740;
    rom_re[76] = -9512;
    rom_re[77] = -10279;
    rom_re[78] = -11039;
    rom_re[79] = -11793;
    rom_re[80] = -12540;
    rom_re[81] = -13279;
    rom_re[82] = -14010;
    rom_re[83] = -14733;
    rom_re[84] = -15447;
    rom_re[85] = -16151;
    rom_re[86] = -16846;
    rom_re[87] = -17531;
    rom_re[88] = -18205;
    rom_re[89] = -18868;
    rom_re[90] = -19520;
    rom_re[91] = -20160;
    rom_re[92] = -20788;
    rom_re[93] = -21403;
    rom_re[94] = -22006;
    rom_re[95] = -22595;
    rom_re[96] = -23170;
    rom_re[97] = -23732;
    rom_re[98] = -24279;
    rom_re[99] = -24812;
    rom_re[100] = -25330;
    rom_re[101] = -25833;
    rom_re[102] = -26320;
    rom_re[103] = -26791;
    rom_re[104] = -27246;
    rom_re[105] = -27684;
    rom_re[106] = -28106;
    rom_re[107] = -28511;
    rom_re[108] = -28899;
    rom_re[109] = -29269;
    rom_re[110] = -29622;
    rom_re[111] = -29957;
    rom_re[112] = -30274;
    rom_re[113] = -30572;
    rom_re[114] = -30853;
    rom_re[115] = -31114;
    rom_re[116] = -31357;
    rom_re[117] = -31581;
    rom_re[118] = -31786;
    rom_re[119] = -31972;
    rom_re[120] = -32138;
    rom_re[121] = -32286;
    rom_re[122] = -32413;
    rom_re[123] = -32522;
    rom_re[124] = -32610;
    rom_re[125] = -32679;
    rom_re[126] = -32729;
    rom_re[127] = -32758;
    rom_im[0] = 0;
    rom_im[1] = -804;
    rom_im[2] = -1608;
    rom_im[3] = -2411;
    rom_im[4] = -3212;
    rom_im[5] = -4011;
    rom_im[6] = -4808;
    rom_im[7] = -5602;
    rom_im[8] = -6393;
    rom_im[9] = -7180;
    rom_im[10] = -7962;
    rom_im[11] = -8740;
    rom_im[12] = -9512;
    rom_im[13] = -10279;
    rom_im[14] = -11039;
    rom_im[15] = -11793;
    rom_im[16] = -12540;
    rom_im[17] = -13279;
    rom_im[18] = -14010;
    rom_im[19] = -14733;
    rom_im[20] = -15447;
    rom_im[21] = -16151;
    rom_im[22] = -16846;
    rom_im[23] = -17531;
    rom_im[24] = -18205;
    rom_im[25] = -18868;
    rom_im[26] = -19520;
    rom_im[27] = -20160;
    rom_im[28] = -20788;
    rom_im[29] = -21403;
    rom_im[30] = -22006;
    rom_im[31] = -22595;
    rom_im[32] = -23170;
    rom_im[33] = -23732;
    rom_im[34] = -24279;
    rom_im[35] = -24812;
    rom_im[36] = -25330;
    rom_im[37] = -25833;
    rom_im[38] = -26320;
    rom_im[39] = -26791;
    rom_im[40] = -27246;
    rom_im[41] = -27684;
    rom_im[42] = -28106;
    rom_im[43] = -28511;
    rom_im[44] = -28899;
    rom_im[45] = -29269;
    rom_im[46] = -29622;
    rom_im[47] = -29957;
    rom_im[48] = -30274;
    rom_im[49] = -30572;
    rom_im[50] = -30853;
    rom_im[51] = -31114;
    rom_im[52] = -31357;
    rom_im[53] = -31581;
    rom_im[54] = -31786;
    rom_im[55] = -31972;
    rom_im[56] = -32138;
    rom_im[57] = -32286;
    rom_im[58] = -32413;
    rom_im[59] = -32522;
    rom_im[60] = -32610;
    rom_im[61] = -32679;
    rom_im[62] = -32729;
    rom_im[63] = -32758;
    rom_im[64] = -32768;
    rom_im[65] = -32758;
    rom_im[66] = -32729;
    rom_im[67] = -32679;
    rom_im[68] = -32610;
    rom_im[69] = -32522;
    rom_im[70] = -32413;
    rom_im[71] = -32286;
    rom_im[72] = -32138;
    rom_im[73] = -31972;
    rom_im[74] = -31786;
    rom_im[75] = -31581;
    rom_im[76] = -31357;
    rom_im[77] = -31114;
    rom_im[78] = -30853;
    rom_im[79] = -30572;
    rom_im[80] = -30274;
    rom_im[81] = -29957;
    rom_im[82] = -29622;
    rom_im[83] = -29269;
    rom_im[84] = -28899;
    rom_im[85] = -28511;
    rom_im[86] = -28106;
    rom_im[87] = -27684;
    rom_im[88] = -27246;
    rom_im[89] = -26791;
    rom_im[90] = -26320;
    rom_im[91] = -25833;
    rom_im[92] = -25330;
    rom_im[93] = -24812;
    rom_im[94] = -24279;
    rom_im[95] = -23732;
    rom_im[96] = -23170;
    rom_im[97] = -22595;
    rom_im[98] = -22006;
    rom_im[99] = -21403;
    rom_im[100] = -20788;
    rom_im[101] = -20160;
    rom_im[102] = -19520;
    rom_im[103] = -18868;
    rom_im[104] = -18205;
    rom_im[105] = -17531;
    rom_im[106] = -16846;
    rom_im[107] = -16151;
    rom_im[108] = -15447;
    rom_im[109] = -14733;
    rom_im[110] = -14010;
    rom_im[111] = -13279;
    rom_im[112] = -12540;
    rom_im[113] = -11793;
    rom_im[114] = -11039;
    rom_im[115] = -10279;
    rom_im[116] = -9512;
    rom_im[117] = -8740;
    rom_im[118] = -7962;
    rom_im[119] = -7180;
    rom_im[120] = -6393;
    rom_im[121] = -5602;
    rom_im[122] = -4808;
    rom_im[123] = -4011;
    rom_im[124] = -3212;
    rom_im[125] = -2411;
    rom_im[126] = -1608;
    rom_im[127] = -804;
  end

  always_comb begin
    re = rom_re[addr];
    im = rom_im[addr];
  end

endmodule
